`timescale 1ns/1ps
module ASYNC_FIFO_tb();
parameter data_width = 8;
  // DUT inputs/outputs

   reg wclk;
   reg wrst_n;
   reg winc;
   reg rclk;
   reg rrst_n;
   reg rinc;
   reg [data_width-1:0] wr_data;
   wire wfull;
   wire rempty;
   wire [data_width-1:0] rd_data;

  // Instantiate DUT
ASYNC_FIFO #(
    .data_width(8),.addr_size(3)
) dut(
    wclk,
    wrst_n,
    winc,
    rclk,
    rrst_n,
    rinc,
    wr_data,
    wfull,
    rempty,
    rd_data
);
  // Clock generation
integer i,j;
parameter reading_clk_freq = 40*10**6;
parameter WRITING_clk_freq = 100*10**6;

parameter reading_clk = 1/(2.0*(reading_clk_freq));
parameter writing_clk = 1/(2.0*(WRITING_clk_freq));

always #12.5 rclk = ~rclk;
always #5    wclk = ~wclk;

initial begin
    $dumpfile("ASYNC_FIFO.vcd");     
    $dumpvars;

    fork
        begin //read
            initialize_r;
            reset_r;
            $display("Start reading 6 bytes...");
                for (j = 0; j < 13; j = j + 1) begin
                    reading(j+1);
                end
                $display("reading is finished");
        
            $stop;

        end
        begin //write
            initialize_w;
            reset_w;
            @(negedge wclk); 
           $display("Start writing 7 bytes...");
                for (i = 0; i < 12; i = i + 1) begin
                    writing(i+1);
                    $display("[%0t] WROTE: %0d", $time, i+1);
                end
          
            $stop;

        end
    join
    #(reading_clk*5);
    $stop;
end
//***********tasks***********//

task reading(input [data_width-1:0] data);
begin
    @(negedge rclk);
    rinc =1;
    @(negedge rclk);
    rinc = 0;
    if (rd_data == data)
            $display("%0t PASS: Expected %0h, Got %0h",$time,data, rd_data);
        else
            $display("%0t FAIL: Expected %0h, Got %0h",$time,data, rd_data);
end
endtask

task writing (input [data_width-1:0] data);
begin
    @(negedge wclk);
    while (wfull) begin
        $display("%0t   FIFO is FULL...", $time);
        @(negedge wclk);
    end
    wr_data = data;
    @(negedge wclk);
    winc = 1;
    @(negedge wclk);
    winc = 0;
end
endtask

task initialize_r;
begin
    rclk = 0;
    rrst_n = 1;
    rinc =0;
end
endtask

task initialize_w;
begin
    wclk = 0;
    wrst_n = 1;
    winc =0;
    wr_data = 8'h00;
    @(negedge wclk);  
end
endtask

task reset_r;
begin
    rrst_n = 1;
    @(negedge rclk);
    rrst_n = 0;
    @(negedge rclk);
    rrst_n = 1;
    @(negedge rclk);

end
endtask
task reset_w;
begin
    wrst_n = 1;
    @(negedge wclk);
    wrst_n = 0;
    @(negedge wclk);
    wrst_n = 1;
    @(negedge wclk);

end
endtask


endmodule